module l2_cache(input clk, input [10:0] address, input l1_miss, output reg hit, output reg miss, output reg [31:0] data_out);
  parameter CACHE_SIZE = 512;
  parameter BLOCK_SIZE = 32;
  parameter NUM_BLOCKS = CACHE_SIZE / BLOCK_SIZE;

  reg valid[NUM_BLOCKS-1:0];
  reg [2:0] tags[NUM_BLOCKS-1:0];
  reg [31:0] data[NUM_BLOCKS-1:0];

  // For a direct-mapped L2 cache with 16 blocks (512/32):
  // Block offset: 5 bits (log2(32) = 5)
  // Index: 4 bits (2^4 = 16 blocks)
  // Tag: 2 bits (11 - 5 - 4 = 2 bits from the address)
  wire [4:0] block_offset = address[4:0];
  wire [3:0] index = address[8:5];
  wire [1:0] tag = address[10:9];

  integer i;
  
  initial begin
    for (i = 0; i < NUM_BLOCKS; i = i + 1) begin
      valid[i] = 0;
    end
  end

  always @(posedge clk) begin
    if (l1_miss) begin
      if (valid[index] && tags[index] == tag) begin
        hit <= 1;
        miss <= 0;
        data_out <= data[index];
        $display("L2 Cache HIT: Address=%h, Index=%h, Tag=%h", address, index, tag);
      end else begin
        hit <= 0;
        miss <= 1;
        data_out <= 0;
        $display("L2 Cache MISS: Address=%h, Index=%h, Tag=%h", address, index, tag);
        // On a miss, we update the cache with data that would come from memory
        // In this simulation, we'll just mark it as valid and update the tag
        valid[index] <= 1;
        tags[index] <= tag;
        data[index] <= 32'hFEEDFACE; // Placeholder data
      end
    end else begin
      hit <= 0;
      miss <= 0;
    end
  end
endmodule
